* cir file corresponding to the equivalent circuit.
* ���� 1
R1 _net1 Input 1.000000 
C1 _net0 _net1 1.000000 
R_C1 _net0 _net1 1.000000 
D1 _net0 0 DMOD_D1 AREA=1.0 Temp=26.85
R_D1 0 _net0 1.000000 
* ���� 2
R2 _net4 Input 1.000000 
C4 0 _net4 1.000000 
R_C2 0 _net4 1.000000 
* ���� 3
R3 _net3 Input 1.000000 
C3 _net2 _net3 1.000000 
R_C3 _net2 _net3 1.000000 
D3 0 _net2 DMOD_D3 AREA=1.0 Temp=26.85
R_D3 0 _net2 1.000000 
.MODEL DMOD_D1 D (Is= 1.000000 N=1.65 Cj0=4e-12 M=0.333 Vj=0.7 Fc=0.5 Rs=0.0686 Tt=5.76e-09 Ikf=0 Kf=0 Af=1 Bv=75 Ibv=1e-06 Xti=3 Eg=1.11 Tcv=0 Trs=0 Ttt1=0 Ttt2=0 Tm1=0 Tm2=0 Tnom=26.85 )
.MODEL DMOD_D3 D (Is= 1.000000 N=1.65 Cj0=4e-12 M=0.333 Vj=0.7 Fc=0.5 Rs=0.0686 Tt=5.76e-09 Ikf=0 Kf=0 Af=1 Bv=75 Ibv=1e-06 Xti=3 Eg=1.11 Tcv=0 Trs=0 Ttt1=0 Ttt2=0 Tm1=0 Tm2=0 Tnom=26.85 )
.END
